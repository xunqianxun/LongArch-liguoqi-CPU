`timescale 1ps/1ps
`include "define.v"

module SnapShortAndRenameTable (
    input        wire                             Clk           ,
    input        wire                             Rest          ,

    //from free list
    input        wire                                                     

    //to free list 

    //from ROB

    //to LSU 用来给违例情况传递最近的CheckPoint

);
    
    reg  []
endmodule