`timescale 1ps/1ps
`include "../define.v"

module AXIbus (
    input
);
    
endmodule