//Computer resource table 计算资源表，可以取消EU计算资源与cluster Issue Queen 握手，直接查询CRT 获取可用计算资源信息
`timescale 1ps/1ps
`include "define.v"

module Crt (
    ports
);
    
endmodule