`timescale 1ps/1ps
`include "../define.v"

module RefTable (
    input       wire                                    Clk              ,
    input       wire                                    Rest             ,
    
);
    
endmodule