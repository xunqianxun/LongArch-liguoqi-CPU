`timescale 1ps/1ps
`include "../define.v"
`include "DecodeOneWay.v"

module Decode (
    input     wire                             Clk           ,
    input     wire                             Rest          ,
    //for ctrl
    input     wire                             DecodeStopS   ,
    input     wire                             DecodeFlashS  ,
    //output    wire                             DecodeReq     ,
    //from InsrQueue
    input     wire                             InInstPort1  ,
    input     wire                             InInstPort2  ,
    input     wire                             InInstPort3  ,
    input     wire                             InInstPort4  ,
    input     wire      [`InstAddrBus]         InInstAddr1   ,
    input     wire      [`InstDateBus]         InInstDate1   ,
    input     wire                             InInstPart1   ,
    input     wire      [`InstAddrBus]         InInstNAdr1   ,
    input     wire      [`InstAddrBus]         InInstAddr2   ,
    input     wire      [`InstDateBus]         InInstDate2   ,
    input     wire                             InInstPart2   ,
    input     wire      [`InstAddrBus]         InInstNAdr2   ,
    input     wire      [`InstAddrBus]         InInstAddr3   ,
    input     wire      [`InstDateBus]         InInstDate3   ,
    input     wire                             InInstPart3   ,
    input     wire      [`InstAddrBus]         InInstNAdr3   ,
    input     wire      [`InstAddrBus]         InInstAddr4   ,
    input     wire      [`InstDateBus]         InInstDate4   ,
    input     wire                             InInstPart4   ,
    input     wire      [`InstAddrBus]         InInstNAdr4   ,
    //input     wire                             QueueEmpty    ,
    //to  distpatch 
    output    wire      [`InstAddrBus]         Inst1Addr     ,
    output    wire      [`MicOperateCode]      Inst1Opcode   ,
    output    wire                             Inst1SinumA   ,
    output    wire      [25:0]                 Inst1SiDate   ,
    output    wire                             Inst1Sr1Abl   ,
    output    wire      [`ArchRegBUs]          Inst1Sr1Num   ,
    output    wire                             Inst1Sr2Abl   ,   
    output    wire      [`ArchRegBUs]          Inst1Sr2Num   ,
    output    wire                             Insr1WriteA   ,
    output    wire                             Inst1Part     , 
    output    wire      [`InstAddrBus]         Inst1Nadr     ,
    output    wire      [`ArchRegBUs]          Inst1WriteN   ,
    output    wire      [`InstAddrBus]         Inst2Addr     ,
    output    wire      [`MicOperateCode]      Inst2Opcode   ,
    output    wire                             Inst2SinumA   ,
    output    wire      [25:0]                 Inst2SiDate   ,
    output    wire                             Inst2Sr1Abl   ,
    output    wire      [`ArchRegBUs]          Inst2Sr1Num   ,
    output    wire                             Inst2Sr2Abl   ,   
    output    wire      [`ArchRegBUs]          Inst2Sr2Num   ,
    output    wire                             Insr2WriteA   ,
    output    wire      [`ArchRegBUs]          Inst2WriteN   ,
    output    wire                             Inst2Part     , 
    output    wire      [`InstAddrBus]         Inst2Nadr     ,
    output    wire      [`InstAddrBus]         Inst3Addr     ,
    output    wire      [`MicOperateCode]      Inst3Opcode   ,
    output    wire                             Inst3SinumA   ,
    output    wire      [25:0]                 Inst3SiDate   ,
    output    wire                             Inst3Sr1Abl   ,
    output    wire      [`ArchRegBUs]          Inst3Sr1Num   ,
    output    wire                             Inst3Sr2Abl   ,   
    output    wire      [`ArchRegBUs]          Inst3Sr2Num   ,
    output    wire                             Insr3WriteA   ,
    output    wire      [`ArchRegBUs]          Inst3WriteN   ,
    output    wire                             Inst3Part     , 
    output    wire      [`InstAddrBus]         Inst3Nadr     ,
    output    wire      [`InstAddrBus]         Inst4Addr     ,
    output    wire      [`MicOperateCode]      Inst4Opcode   ,
    output    wire                             Inst4SinumA   ,
    output    wire      [25:0]                 Inst4SiDate   ,
    output    wire                             Inst4Sr1Abl   ,
    output    wire      [`ArchRegBUs]          Inst4Sr1Num   ,
    output    wire                             Inst4Sr2Abl   ,   
    output    wire      [`ArchRegBUs]          Inst4Sr2Num   ,
    output    wire                             Insr4WriteA   ,
    output    wire      [`ArchRegBUs]          Inst4WriteN   ,
    output    wire                             Inst4Part     , 
    output    wire      [`InstAddrBus]         Inst4Nadr     
);

    DecodeOneWay u1_DecodeOneWay(
        .Clk          ( Clk          ),
        .Rest         ( Rest         ),
        .DecodeStop   ( DecodeStopS  ),
        .DecodeFlash  ( DecodeFlashS ),
        .InInstDate   ( InInstDate1  ),
        .InInstAddr   ( InInstAddr1  ),
        .InInstPart   ( InInstPart1  ),
        .InInstNAdr   ( InInstNAdr1  ),
        .InInstPort   ( InInstPort1  ),
        .InstAddr     ( Inst1Addr    ),
        .InstOpcode   ( Inst1Opcode  ),
        .InstSinumA   ( Inst1SinumA  ),
        .InstSiDate   ( Inst1SiDate  ),
        .InstSr1Abl   ( Inst1Sr1Abl  ),
        .InstSr1Num   ( Inst1Sr1Num  ),
        .InstSr2Abl   ( Inst1Sr2Abl  ),
        .InstSr2Num   ( Inst1Sr2Num  ),
        .InsrWriteA   ( Insr1WriteA  ),
        .InstWriteN   ( Inst1WriteN  ),
        .InstPart     ( Inst1Part    ),
        .InstNadr     ( Inst1Nadr    )
    );

    DecodeOneWay u2_DecodeOneWay(
        .Clk          ( Clk          ),
        .Rest         ( Rest         ),
        .DecodeStop   ( DecodeStopS  ),
        .DecodeFlash  ( DecodeFlashS ),
        .InInstDate   ( InInstDate2  ),
        .InInstAddr   ( InInstAddr2  ),
        .InInstPart   ( InInstPart2  ),
        .InInstNAdr   ( InInstNAdr2  ),
        .InInstPort   ( InInstPort2  ),
        .InstAddr     ( Inst2Addr    ),
        .InstOpcode   ( Inst2Opcode  ),
        .InstSinumA   ( Inst2SinumA  ),
        .InstSiDate   ( Inst2SiDate  ),
        .InstSr1Abl   ( Inst2Sr1Abl  ),
        .InstSr1Num   ( Inst2Sr1Num  ),
        .InstSr2Abl   ( Inst2Sr2Abl  ),
        .InstSr2Num   ( Inst2Sr2Num  ),
        .InsrWriteA   ( Insr2WriteA  ),
        .InstWriteN   ( Inst2WriteN  ),
        .InstPart     ( Inst2Part    ),
        .InstNadr     ( Inst2Nadr    )
    );

    DecodeOneWay u3_DecodeOneWay(
        .Clk          ( Clk          ),
        .Rest         ( Rest         ),
        .DecodeStop   ( DecodeStopS  ),
        .DecodeFlash  ( DecodeFlashS ),
        .InInstDate   ( InInstDate3  ),
        .InInstAddr   ( InInstAddr3  ),
        .InInstPart   ( InInstPart3  ),
        .InInstNAdr   ( InInstNAdr3  ),
        .InInstPort   ( InInstPort3  ),
        .InstAddr     ( Inst3Addr    ),
        .InstOpcode   ( Inst3Opcode  ),
        .InstSinumA   ( Inst3SinumA  ),
        .InstSiDate   ( Inst3SiDate  ),
        .InstSr1Abl   ( Inst3Sr1Abl  ),
        .InstSr1Num   ( Inst3Sr1Num  ),
        .InstSr2Abl   ( Inst3Sr2Abl  ),
        .InstSr2Num   ( Inst3Sr2Num  ),
        .InsrWriteA   ( Insr3WriteA  ),
        .InstWriteN   ( Inst3WriteN  ),
        .InstPart     ( Inst3Part    ),
        .InstNadr     ( Inst3Nadr    )
    );

    DecodeOneWay u4_DecodeOneWay(
        .Clk          ( Clk          ),
        .Rest         ( Rest         ),
        .DecodeStop   ( DecodeStopS  ),
        .DecodeFlash  ( DecodeFlashS ),
        .InInstDate   ( InInstDate4  ),
        .InInstAddr   ( InInstAddr4  ),
        .InInstPart   ( InInstPart4  ),
        .InInstNAdr   ( InInstNAdr4  ),
        .InInstPort   ( InInstPort4  ),
        .InstAddr     ( Inst4Addr    ),
        .InstOpcode   ( Inst4Opcode  ),
        .InstSinumA   ( Inst4SinumA  ),
        .InstSiDate   ( Inst4SiDate  ),
        .InstSr1Abl   ( Inst4Sr1Abl  ),
        .InstSr1Num   ( Inst4Sr1Num  ),
        .InstSr2Abl   ( Inst4Sr2Abl  ),
        .InstSr2Num   ( Inst4Sr2Num  ),
        .InsrWriteA   ( Insr4WriteA  ),
        .InstWriteN   ( Inst4WriteN  ),
        .InstPart     ( Inst4Part    ),
        .InstNadr     ( Inst4Nadr    )
    );



endmodule
