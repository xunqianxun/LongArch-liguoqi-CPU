`timescale 1ps/1ps
`include "define.v"

module ICacheEntry #(
    parameter 
) (
    ports
);
    
endmodule