`ifndef _SOCDEFINE_H_
`define _SOCDEFINE_H_

`define DEBUG_REPORT 1
`define SYNTHESIZE 1

`endif 
