`ifndef _SOCDEFINE_H_
`define _SOCDEFINE_H_
`define LINTCHECK  1  //编写时打开lint工具对代码进行检查


`endif 
