`include "define.v"
module Decode (
    input     wire                             Clk          ,
    input     wire                             Rest         ,

    input     wire     [`InstAddrBus]          InDecodePc   ,
    input     wire     [`TwoInstDateBus]       InDecodeInst ,
    

);
    
endmodule