`timescale 1ps/1ps
`include "define.v"

module PhysicalRegFile (
    input          wire                                 Clk                 ,
    input          wire                                 Rest                ,
    //inst1 dataL read
    input          wire                                 Inst1ReadLAble      ,
    input          wire        [6:0]                    Inst1ReadLAddr      ,
    output         wire        [`DataBus]               PRFDataToTInst1L    ,
    output         wire                                 PRFsuccessToTInst1L ,
    //inst1 dataR read
    input          wire                                 Inst1ReadRAble      ,
    input          wire        [6:0]                    Inst1ReadRAddr      ,
    output         wire        [`DataBus]               PRFDataToTInst1R    ,
    output         wire                                 PRFsuccessToTInst1R ,
    //inst2 dataL read
    input          wire                                 Inst2ReadLAble      ,
    input          wire        [6:0]                    Inst2ReadLAddr      ,
    output         wire        [`DataBus]               PRFDataToTInst2L    ,
    output         wire                                 PRFsuccessToTInst2L ,
    //inst2 dataR read
    input          wire                                 Inst2ReadRAble      ,
    input          wire        [6:0]                    Inst2ReadRAddr      ,
    output         wire        [`DataBus]               PRFDataToTInst2R    ,
    output         wire                                 PRFsuccessToTInst2R ,
    //inst3 dataL read
    input          wire                                 Inst3ReadLAble      ,
    input          wire        [6:0]                    Inst3ReadLAddr      ,
    output         wire        [`DataBus]               PRFDataToTInst3L    ,
    output         wire                                 PRFsuccessToTInst3L ,
    //inst3 dataR read
    input          wire                                 Inst3ReadRAble      ,
    input          wire        [6:0]                    Inst3ReadRAddr      ,
    output         wire        [`DataBus]               PRFDataToTInst3R    ,
    output         wire                                 PRFsuccessToTInst3R ,
    //inst4 dataL read
    input          wire                                 Inst4ReadLAble      ,
    input          wire        [6:0]                    Inst4ReadLAddr      ,
    output         wire        [`DataBus]               PRFDataToTInst4L    ,
    output         wire                                 PRFsuccessToTInst4L ,
    //inst4 dataR read
    input          wire                                 Inst4ReadRAble      ,
    input          wire        [6:0]                    Inst4ReadRAddr      ,
    output         wire        [`DataBus]               PRFDataToTInst4R    ,
    output         wire                                 PRFsuccessToTInst4R ,
    //ALU1 data write 
    input          wire                                 ALU1WriteAble       ,
    input          wire        [6:0]                    ALU1WriteAddr       ,
    input          wire        [`DataBus]               ALU1WriteData       ,
    //ALU2 data write 
    input          wire                                 ALU2WriteAble       ,
    input          wire        [6:0]                    ALU2WriteAddr       ,
    input          wire        [`DataBus]               ALU2WriteData       ,
    //MLU data write 
    input          wire                                 MLUWriteAble        ,
    input          wire        [6:0]                    MLUWriteAddr        ,
    input          wire        [`DataBus]               MLUWriteData        ,
    //DIV data write 
    input          wire                                 DIVWriteAble        ,
    input          wire        [6:0]                    DIVWriteAddr        ,
    input          wire        [`DataBus]               DIVWriteData        ,
    //BRU data write 
    input          wire                                 BRUWriteAble        ,
    input          wire        [6:0]                    BRUWriteAddr        ,
    input          wire        [`DataBus]               BRUWriteData        ,
    //CSRU data write 
    input          wire                                 CSRUWriteAble       ,
    input          wire        [6:0]                    CSRUWriteAddr       ,
    input          wire        [`DataBus]               CSRUWriteData       ,
    //Load data write 
    input          wire                                 LoadWriteAble       ,
    input          wire        [6:0]                    LoadWriteAddr       ,
    input          wire        [`DataBus]               LoadWriteData       ,
    //From ROB relace some physical reg
    input          wire                                 ROBCommit1Able      ,
    input          wire        [6:0]                    ROBCommit1Addr      ,
    input          wire                                 ROBCommit2Able      ,
    input          wire        [6:0]                    ROBCommit2Addr      ,
    input          wire                                 ROBCommit3Able      ,
    input          wire        [6:0]                    ROBCommit3Addr      ,
    input          wire                                 ROBCommit4Able      ,
    input          wire        [6:0]                    ROBCommit4Addr      ,
    // to Arch reg file  and free list
    output         wire                                 PRFwrite1Able       ,
    output         wire        [6:0]                    PRFwrite1Addr       ,
    output         wire        [`DataBus]               PRFwrite1Date       ,
    output         wire                                 PRFwrite2Able       ,
    output         wire        [6:0]                    PRFwrite2Addr       ,
    output         wire        [`DataBus]               PRFwrite2Date       , 
    output         wire                                 PRFwrite3Able       ,
    output         wire        [6:0]                    PRFwrite3Addr       ,
    output         wire        [`DataBus]               PRFwrite3Date       , 
    output         wire                                 PRFwrite4Able       ,
    output         wire        [6:0]                    PRFwrite4Addr       ,
    output         wire        [`DataBus]               PRFwrite4Date       , 

);

    reg  [32+1-1:0] PhysicalReg [0:127] ;
    // integer PRFLoopClean ;
    // always @(posedge Clk) begin
    //     if(!Rest) begin
    //         for (PRFLoopClean = 0;PRFLoopClean < 128 ;PRFLoopClean = PRFLoopClean+1) begin
    //             PhysicalReg[PRFLoopClean] <= 34'd0 ;
    //         end
    //     end
    //     else begin
            
    //     end
    // end
    localparam EMPTY = 1'b0 ;
    localparam FULL  = 1'b1 ;

    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[0] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[0] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[0] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[0] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[0] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[0] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[0] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[0] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[0] <= 33'd0;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[0] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[0] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[0] <= 33'd0;end
    end

    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[1] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd1)) PhysicalReg[1] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd1)) PhysicalReg[1] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd1))  PhysicalReg[1] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd1))  PhysicalReg[1] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd1))  PhysicalReg[1] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd1)) PhysicalReg[1] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd1)) PhysicalReg[1] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd1)) PhysicalReg[1] <= 33'd0;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd1)) PhysicalReg[1] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd1)) PhysicalReg[1] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd1)) PhysicalReg[1] <= 33'd0;end 
    end

    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ; end 
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd2)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd2)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd2))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd2))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd2))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd2)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd2)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd2)) PhysicalReg[2] <= 33'd0;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd2)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd2)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd2)) PhysicalReg[2] <= 33'd0;end
    end 

    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[3] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd3)) PhysicalReg[3] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd3)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end
    end

    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[4] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd4)) PhysicalReg[4] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd4)) PhysicalReg[4] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd4))  PhysicalReg[4] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd4))  PhysicalReg[4] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd4))  PhysicalReg[4] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd4)) PhysicalReg[4] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd4)) PhysicalReg[4] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd4)) PhysicalReg[4] <= 33'd0;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd4)) PhysicalReg[4] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd4)) PhysicalReg[4] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd4)) PhysicalReg[4] <= 33'd0; end
    end

    always @(posedge Clk) begin
        if(!Rest) begin
            PhysicalReg[5] <= 33'd0 ;
        end
        else begin // when read need check write addr 
            if((ALU1WriteAble) && (ALU1WriteAddr == 7'd5)) PhysicalReg[5] <= {ALU1WriteData, FULL} ;
            if((ALU2WriteAble) && (ALU2WriteAddr == 7'd5)) PhysicalReg[5] <= {ALU2WriteData, FULL} ;
            if((MLUWriteAble)  && (MLUWriteAddr == 7'd5))  PhysicalReg[5] <= {MLUWriteData, FULL}  ;
            if((DIVWriteAble)  && (DIVWriteAddr == 7'd5))  PhysicalReg[5] <= {DIVWriteData, FULL}  ;
            if((BRUWriteAble)  && (BRUWriteAddr == 7'd5))  PhysicalReg[5] <= {BRUWriteData, FULL}  ;
            if((CSRUWriteAble) && (CSRUWriteAddr == 7'd5)) PhysicalReg[5] <= {CSRUWriteData, FULL} ;
            if((LoadWriteAble) && (LoadWriteAddr == 7'd5)) PhysicalReg[5] <= {LoadWriteData, FULL} ;
            if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd5)) PhysicalReg[5] <= 33'd0                 ;
            if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd5)) PhysicalReg[5] <= 33'd0                 ;
            if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd5)) PhysicalReg[5] <= 33'd0                 ;
            if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd5)) PhysicalReg[5] <= 33'd0                 ;
        end
    end

    always @(posedge Clk) begin
        if(!Rest) begin
            PhysicalReg[2] <= 33'd0 ;
        end
        else begin // when read need check write addr 
            if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;
            if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;
            if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;
            if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;
            if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;
            if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;
            if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;
            if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0                 ;
            if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0                 ;
            if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0                 ;
            if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0                 ;
        end
    end

    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
        always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    always @(posedge Clk) begin
        if(!Rest) begin PhysicalReg[2] <= 33'd0 ;end
        else begin if((ALU1WriteAble) && (ALU1WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU1WriteData, FULL} ;if((ALU2WriteAble) && (ALU2WriteAddr == 7'd0)) PhysicalReg[2] <= {ALU2WriteData, FULL} ;if((MLUWriteAble)  && (MLUWriteAddr == 7'd0))  PhysicalReg[2] <= {MLUWriteData, FULL}  ;if((DIVWriteAble)  && (DIVWriteAddr == 7'd0))  PhysicalReg[2] <= {DIVWriteData, FULL}  ;if((BRUWriteAble)  && (BRUWriteAddr == 7'd0))  PhysicalReg[2] <= {BRUWriteData, FULL}  ;if((CSRUWriteAble) && (CSRUWriteAddr == 7'd0)) PhysicalReg[2] <= {CSRUWriteData, FULL} ;if((LoadWriteAble) && (LoadWriteAddr == 7'd0)) PhysicalReg[2] <= {LoadWriteData, FULL} ;if((ROBCommit1Able)&& (ROBCommit1Addr== 7'd0)) PhysicalReg[2] <= 33'd0 ;if((ROBCommit2Able)&& (ROBCommit2Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit3Able)&& (ROBCommit3Addr== 7'd0)) PhysicalReg[2] <= 33'd0;if((ROBCommit4Able)&& (ROBCommit4Addr== 7'd0)) PhysicalReg[2] <= 33'd0;end 
    end
    
    
endmodule