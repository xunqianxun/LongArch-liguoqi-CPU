`timescale 1ps/1ps
`include "IPsetting.v"

module CompressCriq (
    input        wire                                       Clk            ,
    input        wire                                       Rest           ,
    
    input        wire         
);
    
endmodule