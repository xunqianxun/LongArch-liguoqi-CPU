`timescale 1ps/1ps
`include "define.v"

module RegRenameTable (
    input         wire                                  Clk               ,
    input         wire                                  Rest              ,


);

    localparam ARF1 = 
    
endmodule