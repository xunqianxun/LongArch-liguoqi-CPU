`timescale 1ps/1ps
`include "../define.v"

module DCacheStage1 (
    input        wire                                 Clk          ,
    input        wire                                 Rest         ,
    //
);
    
endmodule