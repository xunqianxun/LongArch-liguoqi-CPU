`timescale 1ps/1ps
`include "IPsetting.v"

module FifoCtrl(
    input         wire                            Clk           ,
    input         wire                            Rest          ,


);
    
    

endmodule