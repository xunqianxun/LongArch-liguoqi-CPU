`timescale 1ps/1ps
`include "define.v"

module SnapShortAndRenameTable (
    input        wire                             Clk           ,
    input        wire                             Rest          ,

    //input        wire                             
);
    
endmodule