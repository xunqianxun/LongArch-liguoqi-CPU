`timescale 1ps/1ps
`include "../define.v"

module FTQ (
    input       wire                           Clk          ,
    input       wire                           Rest         ,
);
    
endmodule