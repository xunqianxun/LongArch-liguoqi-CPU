`timescale 1ps/1ps
`include "../define.v"

module BusyTable (
    input       wire                                 Clk             ,
    input       wire                                 Rest            ,
    //for ctrl  
    input       wire                                 BusyStop        ,
    input       wire                                 BusyFlash       ,
    //from Issue
    input       wire                                 UnBusyAble1     ,
    input       wire      [`ReNameRegBUs]            UnBusyAddr1     ,    
    input       wire                                 UnBusyAble2     ,
    input       wire      [`ReNameRegBUs]            UnBusyAddr2     ,   
    input       wire                                 UnBusyAble3     ,
    input       wire      [`ReNameRegBUs]            UnBusyAddr3     ,   
    input       wire                                 UnBusyAble4     ,
    input       wire      [`ReNameRegBUs]            UnBusyAddr4     ,                               
    input       wire                                 UnBusyAble5     ,
    input       wire      [`ReNameRegBUs]            UnBusyAddr5     ,   
    input       wire                                 UnBusyAble6     ,
    input       wire      [`ReNameRegBUs]            UnBusyAddr6     ,  
    input       wire                                 UnBusyAble7     ,
    input       wire      [`ReNameRegBUs]            UnBusyAddr7     ,  
    //from RAT
    input       wire                                 BIn1Src1Able     ,
    input       wire     [`ReNameRegBUs]             BIn1Src1Addr     ,
    input       wire                                 BIn1Src2Able     ,
    input       wire     [`ReNameRegBUs]             BIn1Src2Addr     ,
    input       wire                                 BIn1RdAble       ,
    input       wire     [`ReNameRegBUs]             BIn1RdAddr       ,
    input       wire                                 BIn2Src1Able     ,
    input       wire     [`ReNameRegBUs]             BIn2Src1Addr     ,
    input       wire                                 BIn2Src2Able     ,
    input       wire     [`ReNameRegBUs]             BIn2Src2Addr     ,
    input       wire                                 BIn2RdAble       ,
    input       wire     [`ReNameRegBUs]             BIn2RdAddr       ,
    input       wire                                 BIn3Src1Able     ,
    input       wire     [`ReNameRegBUs]             BIn3Src1Addr     ,
    input       wire                                 BIn3Src2Able     ,
    input       wire     [`ReNameRegBUs]             BIn3Src2Addr     ,
    input       wire                                 BIn3RdAble       ,
    input       wire     [`ReNameRegBUs]             BIn3RdAddr       ,
    input       wire                                 BIn4Src1Able     ,
    input       wire     [`ReNameRegBUs]             BIn4Src1Addr     ,
    input       wire                                 BIn4Src2Able     ,
    input       wire     [`ReNameRegBUs]             BIn4Src2Addr     ,
    input       wire                                 BIn4RdAble       ,
    input       wire     [`ReNameRegBUs]             BIn4RdAddr       ,
    //to IssueQueue
    output       wire                                BOut1Src1Able     ,
    output       wire     [`ReNameRegBUs]            BOut1Src1Addr     ,
    output       wire                                BOut1Src2Able     ,
    output       wire     [`ReNameRegBUs]            BOut1Src2Addr     ,
    output       wire                                BOut1RdAble       ,
    output       wire     [`ReNameRegBUs]            BOut1RdAddr       ,
    output       wire                                BOut2Src1Able     ,
    output       wire     [`ReNameRegBUs]            BOut2Src1Addr     ,
    output       wire                                BOut2Src2Able     ,
    output       wire     [`ReNameRegBUs]            BOut2Src2Addr     ,
    output       wire                                BOut2RdAble       ,
    output       wire     [`ReNameRegBUs]            BOut2RdAddr       ,
    output       wire                                BOut3Src1Able     ,
    output       wire     [`ReNameRegBUs]            BOut3Src1Addr     ,
    output       wire                                BOut3Src2Able     ,
    output       wire     [`ReNameRegBUs]            BOut3Src2Addr     ,
    output       wire                                BOut3RdAble       ,
    output       wire     [`ReNameRegBUs]            BOut3RdAddr       ,
    output       wire                                BOut4Src1Able     ,
    output       wire     [`ReNameRegBUs]            BOut4Src1Addr     ,
    output       wire                                BOut4Src2Able     ,
    output       wire     [`ReNameRegBUs]            BOut4Src2Addr     ,
    output       wire                                BOut4RdAble       ,
    output       wire     [`ReNameRegBUs]            BOut4RdAddr       
);

    reg              BusyTableSign  [0:127] 
    
endmodule