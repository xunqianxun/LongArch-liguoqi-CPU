`timescale 1ps/1ps
`include"define.v"

module moduleName #(
    parameter WIDTH_BTB = 32
) (
    input        wire                                   Clk             ,
    input        wire                                   Rest            ,

    input        wire 
);
    
endmodule