`include "define.v"
module IssueQue (
    
);
    
endmodule