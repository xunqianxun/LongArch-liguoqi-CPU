`ifndef TAGEDEFINE_H_
`define TAGEDEFINE_H_

`define TAGEBANNUM  6 
`define GHRWIDE     72
`define BASEDEEP    128
`define T1DEEP      128
`define T2DEEP      128

`endif

